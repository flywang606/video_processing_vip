module test_tb;

`include "pixel_func_unit.v"


endmodule