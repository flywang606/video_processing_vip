
parameter	BINFILE="./../../binary/image_64_64.bin";
'define PIXEL_DEPTH 'd8
'define MEMOEY_SIZE 'h0010_0000 //8MB